// from https://people.ece.cornell.edu/land/courses/eceprojectsland/STUDENTPROJ/2006to2007/dbb26/dbb28_meng_report.pdf (TIA.v)
module objPixelOn(
  input [7:0] pixelNum,
  input [7:0] objPos,
  input [7:0] objMask,
  input [2:0] objSize,
  output      pixelOn
);

  wire [7:0]  objIndex;
  wire [8:0]  objByteIndex;
  wire        objMaskOn, objPosOn;
  reg         objSizeOn;
  reg [2:0]   objMaskSel;

  assign objIndex = pixelNum - objPos - 8'd1;
  assign objByteIndex = 9'b1 << (objIndex[7:3]);

  always @(*) begin
    case (objSize)
      3'd0: objSizeOn = (objByteIndex & 9'b000000001) != 0;
      3'd1: objSizeOn = (objByteIndex & 9'b000000101) != 0;
      3'd2: objSizeOn = (objByteIndex & 9'b000010001) != 0;
      3'd3: objSizeOn = (objByteIndex & 9'b000010101) != 0;
      3'd4: objSizeOn = (objByteIndex & 9'b100000001) != 0;
      3'd5: objSizeOn = (objByteIndex & 9'b000000011) != 0;
      3'd6: objSizeOn = (objByteIndex & 9'b100010001) != 0;
      3'd7: objSizeOn = (objByteIndex & 9'b000001111) != 0;
    endcase
  end

  always @(*) begin
    case (objSize)
      3'd5: objMaskSel = objIndex[3:1];
      3'd7: objMaskSel = objIndex[4:2];
      default: objMaskSel = objIndex[2:0];
    endcase
  end

  assign objMaskOn = objMask[objMaskSel];
  assign objPosOn = (pixelNum > objPos) && ({1'b0, pixelNum} <= {1'b0, objPos} + 9'd72);
  assign pixelOn = objSizeOn && objMaskOn && objPosOn;

endmodule
