module decorder(
  input [7:0]      INSTR,
  output reg [5:0] OP,
  output reg [3:0] ADDR_MODE
);

`include "params.vh"

  always @(*) begin
    case (INSTR)
      8'h00: begin OP = C_OP_BRK; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h01: begin OP = C_OP_ORA; ADDR_MODE = C_ADDR_MODE_INX; end
      8'h05: begin OP = C_OP_ORA; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h06: begin OP = C_OP_ASL; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h08: begin OP = C_OP_PHP; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h09: begin OP = C_OP_ORA; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'h0a: begin OP = C_OP_ASL; ADDR_MODE = C_ADDR_MODE_ACC; end
      8'h0d: begin OP = C_OP_ORA; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h0e: begin OP = C_OP_ASL; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h10: begin OP = C_OP_BPL; ADDR_MODE = C_ADDR_MODE_REL; end
      8'h11: begin OP = C_OP_ORA; ADDR_MODE = C_ADDR_MODE_INY; end
      8'h15: begin OP = C_OP_ORA; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'h16: begin OP = C_OP_ASL; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'h18: begin OP = C_OP_CLC; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h19: begin OP = C_OP_ORA; ADDR_MODE = C_ADDR_MODE_ABY; end
      8'h1a: begin OP = C_OP_INA; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h1d: begin OP = C_OP_ORA; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'h1e: begin OP = C_OP_ASL; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'h20: begin OP = C_OP_JSR; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h21: begin OP = C_OP_AND; ADDR_MODE = C_ADDR_MODE_INX; end
      8'h24: begin OP = C_OP_BIT; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h25: begin OP = C_OP_AND; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h26: begin OP = C_OP_ROL; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h28: begin OP = C_OP_PLP; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h29: begin OP = C_OP_AND; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'h2a: begin OP = C_OP_ROL; ADDR_MODE = C_ADDR_MODE_ACC; end
      8'h2c: begin OP = C_OP_BIT; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h2d: begin OP = C_OP_AND; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h2e: begin OP = C_OP_ROL; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h30: begin OP = C_OP_BMI; ADDR_MODE = C_ADDR_MODE_REL; end
      8'h31: begin OP = C_OP_AND; ADDR_MODE = C_ADDR_MODE_INY; end
      8'h34: begin OP = C_OP_BIT; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'h35: begin OP = C_OP_AND; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'h36: begin OP = C_OP_ROL; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'h38: begin OP = C_OP_SEC; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h39: begin OP = C_OP_AND; ADDR_MODE = C_ADDR_MODE_ABY; end
      8'h3a: begin OP = C_OP_DEA; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h3c: begin OP = C_OP_BIT; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'h3d: begin OP = C_OP_AND; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'h3e: begin OP = C_OP_ROL; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'h40: begin OP = C_OP_RTI; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h41: begin OP = C_OP_EOR; ADDR_MODE = C_ADDR_MODE_INX; end
      8'h45: begin OP = C_OP_EOR; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h46: begin OP = C_OP_LSR; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h48: begin OP = C_OP_PHA; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h49: begin OP = C_OP_EOR; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'h4a: begin OP = C_OP_LSR; ADDR_MODE = C_ADDR_MODE_ACC; end
      8'h4c: begin OP = C_OP_JMP; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h4d: begin OP = C_OP_EOR; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h4e: begin OP = C_OP_LSR; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h50: begin OP = C_OP_BVC; ADDR_MODE = C_ADDR_MODE_REL; end
      8'h51: begin OP = C_OP_EOR; ADDR_MODE = C_ADDR_MODE_INY; end
      8'h55: begin OP = C_OP_EOR; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'h56: begin OP = C_OP_LSR; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'h58: begin OP = C_OP_CLI; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h59: begin OP = C_OP_EOR; ADDR_MODE = C_ADDR_MODE_ABY; end
      8'h5d: begin OP = C_OP_EOR; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'h5e: begin OP = C_OP_LSR; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'h60: begin OP = C_OP_RTS; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h61: begin OP = C_OP_ADC; ADDR_MODE = C_ADDR_MODE_INX; end
      8'h65: begin OP = C_OP_ADC; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h66: begin OP = C_OP_ROR; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h68: begin OP = C_OP_PLA; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h69: begin OP = C_OP_ADC; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'h6a: begin OP = C_OP_ROR; ADDR_MODE = C_ADDR_MODE_ACC; end
      8'h6c: begin OP = C_OP_JMP; ADDR_MODE = C_ADDR_MODE_IND; end
      8'h6d: begin OP = C_OP_ADC; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h6e: begin OP = C_OP_ROR; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h70: begin OP = C_OP_BVS; ADDR_MODE = C_ADDR_MODE_REL; end
      8'h71: begin OP = C_OP_ADC; ADDR_MODE = C_ADDR_MODE_INY; end
      8'h75: begin OP = C_OP_ADC; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'h76: begin OP = C_OP_ROR; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'h78: begin OP = C_OP_SEI; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h79: begin OP = C_OP_ADC; ADDR_MODE = C_ADDR_MODE_ABY; end
      8'h7d: begin OP = C_OP_ADC; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'h7e: begin OP = C_OP_ROR; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'h81: begin OP = C_OP_STA; ADDR_MODE = C_ADDR_MODE_INX; end
      8'h84: begin OP = C_OP_STY; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h85: begin OP = C_OP_STA; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h86: begin OP = C_OP_STX; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'h88: begin OP = C_OP_DEY; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h89: begin OP = C_OP_BIM; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'h8a: begin OP = C_OP_TXA; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h8c: begin OP = C_OP_STY; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h8d: begin OP = C_OP_STA; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h8e: begin OP = C_OP_STX; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'h90: begin OP = C_OP_BCC; ADDR_MODE = C_ADDR_MODE_REL; end
      8'h91: begin OP = C_OP_STA; ADDR_MODE = C_ADDR_MODE_INY; end
      8'h94: begin OP = C_OP_STY; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'h95: begin OP = C_OP_STA; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'h96: begin OP = C_OP_STX; ADDR_MODE = C_ADDR_MODE_ZPY; end
      8'h98: begin OP = C_OP_TYA; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h99: begin OP = C_OP_STA; ADDR_MODE = C_ADDR_MODE_ABY; end
      8'h9a: begin OP = C_OP_TXS; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'h9d: begin OP = C_OP_STA; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'ha0: begin OP = C_OP_LDY; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'ha1: begin OP = C_OP_LDA; ADDR_MODE = C_ADDR_MODE_INX; end
      8'ha2: begin OP = C_OP_LDX; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'ha4: begin OP = C_OP_LDY; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'ha5: begin OP = C_OP_LDA; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'ha6: begin OP = C_OP_LDX; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'ha8: begin OP = C_OP_TAY; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'ha9: begin OP = C_OP_LDA; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'haa: begin OP = C_OP_TAX; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'hac: begin OP = C_OP_LDY; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'had: begin OP = C_OP_LDA; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'hae: begin OP = C_OP_LDX; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'hb0: begin OP = C_OP_BCS; ADDR_MODE = C_ADDR_MODE_REL; end
      8'hb1: begin OP = C_OP_LDA; ADDR_MODE = C_ADDR_MODE_INY; end
      8'hb4: begin OP = C_OP_LDY; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'hb5: begin OP = C_OP_LDA; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'hb6: begin OP = C_OP_LDX; ADDR_MODE = C_ADDR_MODE_ZPY; end
      8'hb8: begin OP = C_OP_CLV; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'hb9: begin OP = C_OP_LDA; ADDR_MODE = C_ADDR_MODE_ABY; end
      8'hba: begin OP = C_OP_TSX; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'hbc: begin OP = C_OP_LDY; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'hbd: begin OP = C_OP_LDA; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'hbe: begin OP = C_OP_LDX; ADDR_MODE = C_ADDR_MODE_ABY; end
      8'hc0: begin OP = C_OP_CPY; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'hc1: begin OP = C_OP_CMP; ADDR_MODE = C_ADDR_MODE_INX; end
      8'hc4: begin OP = C_OP_CPY; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'hc5: begin OP = C_OP_CMP; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'hc6: begin OP = C_OP_DEC; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'hc8: begin OP = C_OP_INY; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'hc9: begin OP = C_OP_CMP; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'hca: begin OP = C_OP_DEX; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'hcc: begin OP = C_OP_CPY; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'hcd: begin OP = C_OP_CMP; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'hce: begin OP = C_OP_DEC; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'hd0: begin OP = C_OP_BNE; ADDR_MODE = C_ADDR_MODE_REL; end
      8'hd1: begin OP = C_OP_CMP; ADDR_MODE = C_ADDR_MODE_INY; end
      8'hd5: begin OP = C_OP_CMP; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'hd6: begin OP = C_OP_DEC; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'hd8: begin OP = C_OP_CLD; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'hd9: begin OP = C_OP_CMP; ADDR_MODE = C_ADDR_MODE_ABY; end
      8'hdd: begin OP = C_OP_CMP; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'hde: begin OP = C_OP_DEC; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'he0: begin OP = C_OP_CPX; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'he1: begin OP = C_OP_SBC; ADDR_MODE = C_ADDR_MODE_INX; end
      8'he4: begin OP = C_OP_CPX; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'he5: begin OP = C_OP_SBC; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'he6: begin OP = C_OP_INC; ADDR_MODE = C_ADDR_MODE_ZPG; end
      8'he8: begin OP = C_OP_INX; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'he9: begin OP = C_OP_SBC; ADDR_MODE = C_ADDR_MODE_IMM; end
      8'hea: begin OP = C_OP_NOP; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'hec: begin OP = C_OP_CPX; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'hed: begin OP = C_OP_SBC; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'hee: begin OP = C_OP_INC; ADDR_MODE = C_ADDR_MODE_ABS; end
      8'hf0: begin OP = C_OP_BEQ; ADDR_MODE = C_ADDR_MODE_REL; end
      8'hf1: begin OP = C_OP_SBC; ADDR_MODE = C_ADDR_MODE_INY; end
      8'hf5: begin OP = C_OP_SBC; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'hf6: begin OP = C_OP_INC; ADDR_MODE = C_ADDR_MODE_ZPX; end
      8'hf8: begin OP = C_OP_SED; ADDR_MODE = C_ADDR_MODE_IMP; end
      8'hf9: begin OP = C_OP_SBC; ADDR_MODE = C_ADDR_MODE_ABY; end
      8'hfd: begin OP = C_OP_SBC; ADDR_MODE = C_ADDR_MODE_ABX; end
      8'hfe: begin OP = C_OP_INC; ADDR_MODE = C_ADDR_MODE_ABX; end
      default: begin OP = 6'hxx; ADDR_MODE = 4'hx; end
   endcase
 end

endmodule
